
package uvm_easy_mam_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    `include "uvm_easy_mam.svh"
endpackage

